// Ripple Carry Adder using Dataflow
module HA(S, C, A, B);       //half adder design
    input A, B;
    output S, C;

    assign S = A ^ B;
    assign C = A & B;
endmodule

module FA(S, C, A, B, Cin);    //full adder design
    input A, B, Cin;
    output S, C;

    assign S = A ^ B ^ Cin;
    assign C = (A & B) | (B & Cin) | (A & Cin);
endmodule

module RCA2(S, Cout, A, B, Cin);   //ripple adder design
    input [3:0] A, B;
    input Cin;
    output [3:0] S;
    output Cout;
    wire [2:0] C;  // Internal carry wires

   
    FA fa0(S[0], C[0], A[0], B[0], Cin);
    FA fa1(S[1], C[1], A[1], B[1], C[0]);
    FA fa2(S[2], C[2], A[2], B[2], C[1]);
    FA fa3(S[3], Cout, A[3], B[3], C[2]);
endmodule

module RCA_tb2();    //test bench of ripple carry adder
    reg [3:0] A, B;
    reg Cin;
    wire [3:0] S;
    wire Cout;

    RCA rr(S, Cout, A, B, Cin);
    
    initial begin
        A = 4'b0000; B = 4'b0001; Cin = 1'b0;
        #20;
        A = 4'b0101; B = 4'b0011; Cin = 1'b0;
    end
    
    initial 
        $monitor("A=%b B=%b Sum=%b Cout=%b", A, B, S, Cout);
endmodule
